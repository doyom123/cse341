module cla();


endmodule



module alu();

endmodule